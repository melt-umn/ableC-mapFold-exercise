grammar edu:umn:cs:melt:exts:ableC:mapFold;

exports edu:umn:cs:melt:exts:ableC:mapFold:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:mapFold:concretesyntax;

